-- John Taylor, Preeti Chitre, Joel Montes de Oca, Fabian Rosadi
-- Cal Poly Pomona, Spring 2001

-- ALU entity
-- OPERATION  Name           Function
-- 0000       AND            Z <= A and B
-- 0001       OR             Z <= A or B
-- 0010       XOR            Z <= A xor B
-- 0011       NOT (invert)   Z <= not A
-- 0100       ADD            Z <= A + B
-- 0101       SUBtract       Z <= A - B
-- 0110       ROtate Left    Z <= A<14:0> & A<15>
-- 0111       Rotate Right   Z <= A<0> & A<15:1>
-- 1000       SHift Left     Z <= A<14:0> & B<0>
-- 1001       Shift Right    Z <= B<0> & A<15:1>

-- Flags ZERO, CARRY, OVERFLOW, NEGATIVE are generated as appropriate.
-- To generate a CARRY for addition and subtraction, the operands are
-- expanded to 17 bits, where the 17th bit represents the carry.
-- OVERFLOW is generated by XORing the last carry bit with the previous
-- two carries.

-- All shifts and rotates are shifted or rotated one bit.  The bit being
-- shifted out or rotated goes to the CARRY flag.  The LSB of signal B
-- becomes the bit being shifted in for the shift operations.

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

entity ALU is
   port (A, B: in STD_LOGIC_VECTOR (15 downto 0);
         OPERATION: in STD_LOGIC_VECTOR (3 downto 0);
         Z: out STD_LOGIC_VECTOR (15 downto 0);
         ZERO, CARRY, OVERFLOW, NEGATIVE: out STD_LOGIC
   );
end entity;

architecture inside of ALU is

-- Signal to receive the output of the ALU before going to the output port
signal ALU_OUT: STD_LOGIC_VECTOR (15 downto 0);

-- Output of the adder/subtractor
signal SUM: STD_LOGIC_VECTOR (16 downto 0);

constant ALU_AND: STD_LOGIC_VECTOR (3 downto 0) := "0000";
constant ALU_OR : STD_LOGIC_VECTOR (3 downto 0) := "0001";
constant ALU_XOR: STD_LOGIC_VECTOR (3 downto 0) := "0010";
constant ALU_NOT: STD_LOGIC_VECTOR (3 downto 0) := "0011";
constant ALU_ADD: STD_LOGIC_VECTOR (3 downto 0) := "0100";
constant ALU_SUB: STD_LOGIC_VECTOR (3 downto 0) := "0101";
constant ALU_ROL: STD_LOGIC_VECTOR (3 downto 0) := "0110";
constant ALU_ROR: STD_LOGIC_VECTOR (3 downto 0) := "0111";
constant ALU_SHL: STD_LOGIC_VECTOR (3 downto 0) := "1000";
constant ALU_SHR: STD_LOGIC_VECTOR (3 downto 0) := "1001";

begin
   process (OPERATION, A, B, ALU_OUT, SUM)
   begin
      case OPERATION is
         -- ADD operation
         when ALU_ADD =>
            SUM <= (('0' & A) + ('0' & B));
            ALU_OUT <= SUM(15 downto 0);
            CARRY <= SUM(16);
            OVERFLOW <= A(14) xor B(14) xor SUM(14) xor SUM(16);

         -- SUB operation
         when ALU_SUB =>
            SUM <= (('0' & A) + ('0' & (not B))) + '1';
            ALU_OUT <= SUM(15 downto 0);
            CARRY <= SUM(16);
            OVERFLOW <= A(14) xor (not B(14)) xor SUM(14) xor SUM(16);

         -- AND operation
         when ALU_AND =>
            SUM <= "-----------------";
            ALU_OUT <= A and B;
            OVERFLOW <= '0';
            CARRY <= '0';

         -- OR operation
         when ALU_OR =>
            SUM <= "-----------------";
            ALU_OUT <= A or B;
            OVERFLOW <= '0';
            CARRY <= '0';

         -- XOR operation
         when ALU_XOR =>
            SUM <= "-----------------";
            ALU_OUT <= A xor B;
            OVERFLOW <= '0';
            CARRY <= '0';

         -- NOT operation
         when ALU_NOT =>
            SUM <= "-----------------";
            ALU_OUT <= not A;
            OVERFLOW <= '0';
            CARRY <= '0';

         when ALU_ROL =>
            SUM <= "-----------------";
            ALU_OUT <= A(14 downto 0) & A(15);
            OVERFLOW <= '0';
            CARRY <= A(15);

         when ALU_ROR =>
            SUM <= "-----------------";
            ALU_OUT <= A(0) & A(15 downto 1);
            OVERFLOW <= '0';
            CARRY <= A(0);

         when ALU_SHL =>
            SUM <= "-----------------";
            ALU_OUT <= A(14 downto 0) & B(0);
            OVERFLOW <= '0';
            CARRY <= A(15);

         when ALU_SHR =>
            SUM <= "-----------------";
            ALU_OUT <= B(0) & A(15 downto 1);
            OVERFLOW <= '0';
            CARRY <= A(0);

         -- others
         when others =>
            SUM <= "-----------------";
            ALU_OUT <= "----------------";
            OVERFLOW <= '-';
            CARRY <= '-';
      end case;

      -- Determine ZERO flag
      if ALU_OUT(15 downto 0) = "0000000000000000" then
         ZERO <= '1';
      else
         ZERO <= '0';
      end if;
   end process;

   NEGATIVE <= ALU_OUT(15);

   Z <= ALU_OUT(15 downto 0);
end architecture;


